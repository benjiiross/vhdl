library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity buffered_alu_testbench is
end buffered_alu_testbench;

architecture testbench of buffered_alu_testbench is
end architecture testbench;